library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity tb_TOP is

end tb_TOP;

architecture ARCH_1 of tb_TOP is

	

	begin

end ARCH_1;

