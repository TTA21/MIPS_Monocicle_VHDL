library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity MUX_2_5_5 is

port(

	i_INPUT_1_5    :   in std_logic_vector(4 downto 0);
    i_INPUT_2_5    :   in std_logic_vector(4 downto 0);
    i_SEL_2         :   in std_logic;
    o_OUT_5        :   out std_logic_vector(4 downto 0)

);

end MUX_2_5_5;

architecture ARCH_1 of MUX_2_5_5 is

	begin

    o_OUT_5    <=  i_INPUT_1_5 when i_SEL_2 = '0' else i_INPUT_2_5;
	
end ARCH_1;